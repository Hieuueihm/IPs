module key_expansion(
	input clk,
	input rst_n,

	input [127:0] key_i,
	input valid_i,


	);

endmodule