module aes_controller(
	input clk,
	input rst_n,
	input start_i,

	);


	localparam 
	


endmodule